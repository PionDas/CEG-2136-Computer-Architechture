library verilog;
use verilog.vl_types.all;
entity lab3top_vlg_vec_tst is
end lab3top_vlg_vec_tst;

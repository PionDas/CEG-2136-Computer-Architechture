library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity input_generator_low_freq is
port(clk: in std_logic;
     code0: in std_logic;
	  code1: in std_logic;
	  code2: in std_logic;
     S0: out std_logic;
	  S1: out std_logic;
	  S2: out std_logic;
	  S3: out std_logic;
	  A0: out std_logic;
	  A1: out std_logic;
	  A2: out std_logic;
	  A3: out std_logic;
	  B0: out std_logic;
	  B1: out std_logic;
	  B2: out std_logic;
	  B3: out std_logic
     );
end input_generator_low_freq;

architecture behavioral of input_generator_low_freq is
type states is (state0,state1,state2,state3,state4,state5,state6,state7,state8,state9,state10,state11,state12,state13,state14,state15);
signal pr_state, nx_state: states; 
signal my_clk: std_logic;
begin
process(clk)
variable count: integer range 0 to 63000000;
begin
if (clk'event and clk='0')then
	if (count=63000000) then
		my_clk <= not my_clk;
		count:=0;
	else
		count:=count+1;
	end if;
end if;
end process;

process(my_clk)
begin
if (my_clk'event and my_clk='0') then
	pr_state <= nx_state;
end if;
end process;

process(pr_state)
variable reset: std_logic := '1';
begin
if (reset='1') then
	nx_state <= state0;
	reset:='0';
else
	if code0='0' and code1='0' and code2='0' then
		case(pr_state) is
			when state0 => 
				nx_state <=state1;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state1 =>
				nx_state <=state2;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state2 =>
				nx_state <=state3;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state3 =>
				nx_state <=state4;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state4 =>
				nx_state <=state5;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state5 =>
				nx_state <=state6;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state6 =>
				nx_state <=state7;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state7 =>
				nx_state <=state8;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state8 =>
				nx_state <=state9;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state9 =>
				nx_state <=state10;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state10 =>
				nx_state <=state11;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state11 =>
				nx_state <=state12;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state12 =>
				nx_state <=state13;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state13 =>
				nx_state <=state14;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state14 =>
				nx_state <=state15;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			when state15 =>
				nx_state <=state0;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='1';
				B2 <='0';
				B3 <='0';
			end case;
	elsif code0='1' and code1='0' and code2='0' then
		case(pr_state) is
			when state0 => 
				nx_state <=state1;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state1 =>
				nx_state <=state2;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state2 =>
				nx_state <=state3;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state3 =>
				nx_state <=state4;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state4 =>
				nx_state <=state5;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state5 =>
				nx_state <=state6;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state6 =>
				nx_state <=state7;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state7 =>
				nx_state <=state8;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state8 =>
				nx_state <=state9;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state9 =>
				nx_state <=state10;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state10 =>
				nx_state <=state11;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state11 =>
				nx_state <=state12;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state12 =>
				nx_state <=state13;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state13 =>
				nx_state <=state14;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state14 =>
				nx_state <=state15;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			when state15 =>
				nx_state <=state0;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='1';
				A3 <='0';
				B0 <='1';
				B1 <='0';
				B2 <='1';
				B3 <='0';
			end case;
	elsif code0='0' and code1='1' and code2='0' then
		case(pr_state) is
			when state0 => 
				nx_state <=state1;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state1 =>
				nx_state <=state2;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state2 =>
				nx_state <=state3;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state3 =>
				nx_state <=state4;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state4 =>
				nx_state <=state5;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state5 =>
				nx_state <=state6;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state6 =>
				nx_state <=state7;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state7 =>
				nx_state <=state8;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state8 =>
				nx_state <=state9;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state9 =>
				nx_state <=state10;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state10 =>
				nx_state <=state11;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state11 =>
				nx_state <=state12;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state12 =>
				nx_state <=state13;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state13 =>
				nx_state <=state14;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state14 =>
				nx_state <=state15;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			when state15 =>
				nx_state <=state0;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='1';
				A2 <='0';
				A3 <='1';
				B0 <='0';
				B1 <='0';
				B2 <='1';
				B3 <='1';
			end case;
	elsif code0='1' and code1='1' and code2='0' then
		case(pr_state) is
			when state0 => 
				nx_state <=state1;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state1 =>
				nx_state <=state2;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state2 =>
				nx_state <=state3;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';	
			when state3 =>
				nx_state <=state4;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state4 =>
				nx_state <=state5;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state5 =>
				nx_state <=state6;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state6 =>
				nx_state <=state7;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state7 =>
				nx_state <=state8;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state8 =>
				nx_state <=state9;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state9 =>
				nx_state <=state10;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state10 =>
				nx_state <=state11;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state11 =>
				nx_state <=state12;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state12 =>
				nx_state <=state13;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state13 =>
				nx_state <=state14;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state14 =>
				nx_state <=state15;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			when state15 =>
				nx_state <=state0;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='0';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='1';
				B2 <='1';
				B3 <='0';
			end case;
	elsif code0='0' and code1='0' and code2='1' then
		case(pr_state) is
			when state0 => 
				nx_state <=state1;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state1 =>
				nx_state <=state2;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state2 =>
				nx_state <=state3;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state3 =>
				nx_state <=state4;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state4 =>
				nx_state <=state5;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state5 =>
				nx_state <=state6;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state6 =>
				nx_state <=state7;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state7 =>
				nx_state <=state8;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='0';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state8 =>
				nx_state <=state9;
				S0 <='0';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state9 =>
				nx_state <=state10;
				S0 <='1';
				S1 <='0';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state10 =>
				nx_state <=state11;
				S0 <='0';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state11 =>
				nx_state <=state12;
				S0 <='1';
				S1 <='1';
				S2 <='0';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state12 =>
				nx_state <=state13;
				S0 <='0';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state13 =>
				nx_state <=state14;
				S0 <='1';
				S1 <='0';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state14 =>
				nx_state <=state15;
				S0 <='0';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			when state15 =>
				nx_state <=state0;
				S0 <='1';
				S1 <='1';
				S2 <='1';
				S3 <='1';
				A0 <='1';
				A1 <='0';
				A2 <='1';
				A3 <='1';
				B0 <='1';
				B1 <='0';
				B2 <='0';
				B3 <='1';
			end case;
	else 
		S0 <='1';
		S1 <='1';
		S2 <='1';
		S3 <='1';
		A0 <='1';
		A1 <='1';
		A2 <='1';
		A3 <='1';
		B0 <='1';
		B1 <='1';
		B2 <='1';
		B3 <='1';		
	end if;
end if;
end process;

end behavioral;

library verilog;
use verilog.vl_types.all;
entity lab3controller_vlg_vec_tst is
end lab3controller_vlg_vec_tst;
